library verilog;
use verilog.vl_types.all;
entity TestTournamentPredictor is
end TestTournamentPredictor;
