library verilog;
use verilog.vl_types.all;
entity TestGSharePredictor is
end TestGSharePredictor;
