library verilog;
use verilog.vl_types.all;
entity TestPSharePredictor is
end TestPSharePredictor;
